module simple_adder_example (
    input  logic [7:0] a,         // Перше 8-бітне число
    input  logic [7:0] b,         // Друге 8-бітне число
    output logic [7:0] sum_out,   // 8-бітна сума
    output logic       carry_out  // Біт переносу (overflow)
);

    // Оголошуємо проміжний сигнал temp_sum, який має на 1 біт більше,
    // щоб зберігати результат додавання, включаючи можливий перенос.
    // WIDTH (8) + 1 = 9 біт
    logic [8:0] temp_sum;

    // Використовуємо 'always_comb' для комбінаційної логіки.
    // Цей блок буде виконуватись щоразу, коли змінюється 'a' або 'b'.
    always_comb begin
        // Конкатенація '{1'b0, a}' додає нульовий біт до старшого розряду 'a'.
        // Це робиться для того, щоб SystemVerilog розглядав 'a' і 'b' як 9-бітні числа
        // під час додавання, дозволяючи зберегти можливий перенос.
        // Результат додавання зберігається у 9-бітному 'temp_sum'.
        temp_sum = {1'b0, a} + {1'b0, b};
    end

    // Присвоюємо молодші 8 бітів temp_sum до sum_out.
    assign sum_out = temp_sum[7:0];

    // Присвоюємо найстарший біт temp_sum (біт переносу) до carry_out.
    assign carry_out = temp_sum[8];

endmodule